module CMSSbox ( in_1, in_2, i_clk, i_r, out_1, out_2 );
(* SILVER="[3:0]_0" *)  input [3:0] in_1;
(* SILVER="[3:0]_1" *)  input [3:0] in_2;
(* SILVER="refresh" *)  input [11:0] i_r;
(* SILVER="[3:0]_0" *)  output [3:0] out_1;
(* SILVER="[3:0]_1" *)  output [3:0] out_2;
(* SILVER="clock" *)  input i_clk;
